module test;
  
  reg clk,rst;
  wire[2:0]count;
  
  counter dut(clk,rst,count);
  
  initial begin
    clk = 0;
    rst = 1;
    #13 rst = 0;
    #1000 $finish;
  end
  
  always #5 clk =~clk;
  
  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0,clk,rst,count);
  end
  
endmodule
